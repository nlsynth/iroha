module mod_comb(clk, rst_n, arg_0, ret_0);
   input clk;
   input rst_n;
   input [31:0] arg_0;
   output [31:0] ret_0;

   assign ret_0 = arg_0;

endmodule // mod_comb
