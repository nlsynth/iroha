module mod_hello(clk, rst);
   input clk;
   input rst;
endmodule
